`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:42:31 02/01/2019 
// Design Name: 
// Module Name:    ANDER_4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ANDER_4(input [3:0]A,input [3:0]B,output [3:0]Y);
	assign Y=A & B;
endmodule
